`include "test.v"
`include "apb_slave"
